`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/04/2022 01:55:12 PM
// Design Name: 
// Module Name: mainTestbench
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module mainTestbench();
    reg b1 = 0, b2 = 0, b3 = 0, b4 = 0, b5 = 0, b6 = 0, b7 = 0, b8 = 0, b9 = 0; 
    reg clk,rst; 
    wire [0:6] seg; 
    wire [3:0] ano; 
        
    main M(clk, b1, b2, b3, b4, b5, b6, b7, b8, b9, rst, seg, ano);
    
    initial begin 
        clk = 1; 
        forever #5 clk = ~clk;
     end
             
    integer i;
    integer j;
    integer k;
     
    initial begin
        rst = 1;
        #20000000
        rst = 0;
        
       
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            b1 = 1;
            b2 = 1;
            b3 = 1;
            b4 = 1;
            #100
            b1 = 0;
            b2 = 0;
            b3 = 0;
            b4 = 0;
            #100
            
       #20000000
        b7 = 1;
        #20000000
        b7 = 0; 
        #20
        b5 = 1; 
        #20000000
        b5 = 0;
        #20
        b6 = 1; 
        #20000000
        b6 = 0; 
        #20
        b8 = 1; 
        #20000000
        b8 = 0;
        #20
        b9 = 1; 
        #20000000
        b9 = 0; 
        
        b4=1;
        #100
        b4=0;
        #100
        b4=1;
        #100
        b4=0;
        #100
        b4=1;
        #100
        b4=0;
        #100
         b4=1;
        #100
        b4=0;
        #100
        b4=1;
        #100
        b4=0;
        #100
        b4=1;
        #100
        b4=0;
        #100
         b4=1;
        #100
        b4=0;
        #100
        b4=1;
        #100
        b4=0;
        #100
        b4=1;
        #100
        b4=0;
        
        #20000000
        b6 = 1; 
        #20000000
        b6 = 0; 
        #20
        b8 = 1; 
        #20000000
        b8 = 0;
        #20
        b9 = 1;
        #20000000
        b9=0;
        
        b1=1;
        #100
        b1=0;
        #100
        b1=1;
        #100
        b1=0;
        #100
        b1=1;
        #100
        b1=0;
        #100
        b1=1;
        #100
        b1=0;
         
        b2=1;
        #100
        b2=0;
        #100
        b2=1;
        #100
        b2=0;
        #100
        b2=1;
        #100
        b2=0;
        
        
          #20000000
        b6 = 1; 
        #20000000
        b6 = 0; 
        #20
        b8 = 1; 
        #20000000
        b8 = 0;
        #20
        b7 = 1;
        #20000000
        b7 = 0; 
        #20
        b9 = 1;
        #200
        b9=0;
        
        b4=1;
        b3=1;
        #100
        b4=0;
        b3=0;
        #100
        b4=1;
        b3=1;
        #100
        b4=0;
        b3=0;
        
        #20000000
        b8=1;
        
    end   
        
    
    
endmodule

